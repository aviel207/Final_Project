///////////////////////////////////
// Verilog testbench
///////////////////////////////////

`timescale	1ns/1ps

module tb_top
(
);
reg  tb_clk, tb_reset;
reg  button_tx;
reg  tb_RxD;
wire tb_done_M;
wire tb_done_d;
wire tb_done_K;
wire tb_done_L;
wire tb_done_r;
wire tb_done_keylen;
wire tb_done_padding;
wire tb_done_rx;
wire tb_TxD;

initial begin
//  $display ("time\t\t  clk reset	 btn 	 rx 	 tx   ");
//  $monitor ("%8g\t\t%b   %b    %b	%b	%b", 
//	  $time, tb_clk, tb_reset, button_tx , tb_RxD , tb_TxD);	        	
  tb_clk             = 1; 
  tb_reset           = 1;
  button_tx 		 = 0;
  #700   tb_reset    = 0;
  
// message arrival
  #0	    tb_RxD   = 1;
  
  //1: "11" - 11
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //2: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //3: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //4: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //5: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //6: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //7: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //8: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //9: "22" - 12
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //10: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //11: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //12: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //13: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //14: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //15 "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //16: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //17: "33" - 13  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //18: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //19: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //20: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //21: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //22: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //23: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //24: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //25: "44" - 14  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //26: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //27: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //28: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //29: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //30 "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //31: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //32: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //33: "55" - 15  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //34: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //35: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //36: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //37: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //38: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //39: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //40: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //41: "66" - 16  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //42: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //43: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //44: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //45: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //46: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //47: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //48: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //49: "77" - 17  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //50: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //51: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //52: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //53: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //54: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //55: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //56: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //57: "11" - 21
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //58: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //59: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //60: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //61: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //62: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //63: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //64: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //65: "22" - 22
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //66: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //67: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //68: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //69: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //70: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //71: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //72: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //73: "33" - 23  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //74: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //75: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //76: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //77: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //78: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //79: "22" 
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //80: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //81: "44" - 24 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //82: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //83: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //84: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //85: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //86: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //87: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //88: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //89: "55" - 25  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //90: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //91: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //92: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //93: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //94: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //95: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //96: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //97: "66" - 26  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //98: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //99: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //100: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //101: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //102: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //103: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //104: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //105: "77" - 27  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //106: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //107: "22" 
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //108: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //109: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //110: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //111: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //112: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //113: "11" - 31
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //114: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //115: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //116: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //117: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //118: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //119: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //120: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //121: "22" - 32
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //122: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //123: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //124: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //125: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //126: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //127: "11" 
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //128: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //129: "33" - 33 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //130: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //131: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //132: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //133: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //134: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //135: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //136: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //137: "44" - 34  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //138: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //139: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //140: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //141: "11" - 11
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //142: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //143: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //144: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //145: "55" - 35  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //146: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //147: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //148: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //149: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //150: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //151: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //152: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //153: "66" - 36  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //154: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //155: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //156: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //157: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //158: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //159: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //160: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //161: "77" - 37  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //162: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //163: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //164: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //165: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //166: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //167: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //168: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //169: "11" - 41
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //170: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //171: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //172: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //173: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //174: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //175: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //176: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //177: "22" - 42
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //178: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //179: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //180: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //181: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //182: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //183: "11" 
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //184: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //185: "33" - 43  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //186: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //187: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //188: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //189: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //190: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //191: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //192: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //193: "44" - 44  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //194: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //195: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //196: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //197: "11" - 11
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //198: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //199: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //200: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //201: "55" - 45
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //202: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //203: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //204: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //205: "22" 
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //206: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //207: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //208: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //209: "66"  - 46 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //210: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //211: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //212: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //213: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //214: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //215: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //216: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //217: "77" - 47  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //218: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //219: "22" 
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //220: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //221: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //222: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //223: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //224: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //225: "11" - 51
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //226: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //227: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //228: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //229: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //230: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //231: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //232: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //233: "22" - 52
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //234: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //235: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //236: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //237: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //238: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //239: "11" - 11
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //240: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //241: "33" - 53  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //242: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //243: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //244: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //245: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //246: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //247: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //248: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //249:"44" - 54  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //250: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //251: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //252: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //253: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //254: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //255: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //256: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //257: "55" - 55  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //258: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //259: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //260: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //261: "22" 
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //262: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //263: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //264: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //265: "66" - 56 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //266: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //267: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //268: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //269: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //270: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //271: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //272: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //273: "77" - 57  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //274: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //275: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //276: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //277: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //278: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //279: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //280: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //281: "11" - 61
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //282: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //283: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //284: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //285: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //286: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //287: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //288: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //289: "22" - 62
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //290: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //291: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //292: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //293: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //294: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //295: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //296: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //297: "33" - 63  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //298: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //299: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //300: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //301: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //302: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //303: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //304: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //305: "44" - 64  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //306: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //307 :"66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //308: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //309: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //310: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //311: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //312: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //313: "55" - 65  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //314: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //315: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //316: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //317: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //318: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //319: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //320: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //321: "66" - 66  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //322: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //323: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //324: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //325: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //326: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //327: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //328: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //329: "77" - 67  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //330: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //331: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //332: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //333: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //334: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //335: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //336: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //337: "11" - 71
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //338: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //339: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //340: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //341: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //342: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //343: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //344: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //345: "22" - 72
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //346: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //347: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //348: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //349: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //350: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //351: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //352: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //353: "33" - 73  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //354: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //355: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //356: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //357: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //358: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //359: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //360: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //361: "44" - 74  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //362: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //363: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //364: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //365: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //366: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //367: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //368: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //369: "55" - 75  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //370: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //371: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //372: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //373: "22" - 12
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //374: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //375: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //376: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //377: "66" - 76  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //378: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //379: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //380: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //381: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //382: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //383: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //384: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //385: "77" - 77  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //386: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //387: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //388: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //389: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //390: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //391: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //392: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //393: "11" - 81
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //394: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //395: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //396: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //397: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //398: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //399: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //400: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //401: "22" - 82
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //402: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //403: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //404: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //405: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //406: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //407: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //408: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //409: "33" - 83  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //410: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //411: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //412: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //413: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //414: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //415: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //416: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //417: "44" - 84  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //418: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //419: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //420: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //421: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //422: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //423: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //424: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //425: "55" - 85  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //426: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //427: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //428: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //429: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //430: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //431: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //432: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //433: "66" - 86  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //434: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //435: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //436: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //437: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //438: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //439: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //440: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //441: "77" - 87  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //442: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //443: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //444: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //445: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //446: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //447: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //448: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
   //449: "11" - 91
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //450: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //451: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //452: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //453: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //454: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //455: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //456: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //457: "22" - 92
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //458: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //459: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //460: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //461: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //462: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //463: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //464: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //465: "33" - 93  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //466: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //467: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //468: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //469: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //470: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //471: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //472: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //473: "44" - 94  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //474: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //475: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //476: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //477: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //478: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //479: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //480: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //481: "55" - 95  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //482: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //483: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //484: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //485: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //486: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //487: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //488: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //489: "66" - 96  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //490: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //491: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //492: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //493: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //494: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //495: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //496: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //497: "77" - 97  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //498: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //499: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //500: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //501: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //502: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //503: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //504: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //505: "11" - 101
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //506: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //507: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //508: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //509: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //510: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //511: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //512: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //513: "22" - 102
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //514: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //515: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //516: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //517: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //518: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //519: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //520: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //521: "33" - 103  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //522: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //523: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //524: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //525: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //526: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //527: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //528: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //529: "44" - 104  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //530: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //531: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //532: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //533: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //534: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //535: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //536: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //537: "55" - 105  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //538: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //539: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //540: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //541: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //542: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //543: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //544: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //545: "66" - 106  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //546: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //547: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //548: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //549: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //550: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //551: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //552: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //553: "77" - 107  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //554: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //555: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //556: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //557: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //558: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //559: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //560: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //561: "11" - 111
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //562: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //563: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //564: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //565: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //566: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //567: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //568: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //569: "22" - 112
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //570: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //571: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //572: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //573: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //574: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //575: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //576: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //577: "33" - 113  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //578: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //579: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //580: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //581: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //582: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //583: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //584: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //585: "44" - 114  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //586: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //587: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //588: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //589: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //590: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //591: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //592:"44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //593: "55" - 115  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //594: "66"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //595: "77"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //596: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;  
  
  //597: "22"
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //598: "33"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //599: "44"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //600: "55"  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 

 //601 padding zeros
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //602 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //603 padding zeros
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //604 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //605 padding zeros
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 

 //606 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //607 padding zeros
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //608 padding zeros
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //609 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //610 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 

 //611 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //612 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //613 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //614 padding zeros
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //615 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 

 //616 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //617 padding zeros
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //618 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //619 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //620 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //621 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //622 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //623 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //624 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //625 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 

 //626 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //627 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //628 padding zeros 38
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //629 padding zeros 39
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //630 padding zeros 40
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //631 padding zeros 41
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //632 padding zeros 42
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //633 padding zeros 43
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //634 padding zeros 44
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //635 padding zeros 45
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 

 //636 padding zeros 46
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //637 padding zeros 47
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //638 padding zeros 48
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //639 padding zeros 49
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //640 padding zeros 50
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //641 padding zeros 51
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //642 padding zeros 52
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //643 padding zeros 53
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //644 padding zeros 54
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //645 padding zeros 55
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 

 //646 padding zeros 56
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //647 padding zeros 57
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //648 padding zeros 58
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //649 padding zeros 59
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //650 padding zeros 60
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //651 padding zeros 61
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //652 padding zeros 62
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //653 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

 //654 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

 //655 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //656 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //657 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //658 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //659 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

 //660 padding zeros 60
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //661 padding zeros 61
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //662 padding zeros 62
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //663 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

 //664 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

 //665 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //666 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //667 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //668 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //669 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //670 padding zeros 60
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //671 padding zeros 61
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //672 padding zeros 62
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //673 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

 //674 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

 //675 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //676 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //677 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //678 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //679 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //680 padding zeros 60
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //681 padding zeros 61
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //682 padding zeros 62
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //683 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

 //684 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

 //685 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //686 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //687 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //688 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //689 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  //690 padding zeros 60
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //691 padding zeros 61
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //692 padding zeros 62
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //693 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

 //694 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

 //695 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //696 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //697 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //698 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //699 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

 //700 padding zeros  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 

 //701 padding zeros
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //702 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //703 padding zeros
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //704 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //705 padding zeros
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 

 //706 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //707 padding zeros
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //708 padding zeros
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //709 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //710 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 

 //711 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //712 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //713 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //714 padding zeros
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //715 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 

 //716 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //717 padding zeros
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //718 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //719 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //720 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //721 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //722 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //723 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //724 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //725 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 

 //726 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //727 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //728 padding zeros 38
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //729 padding zeros 39
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //730 padding zeros 40
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //731 padding zeros 41
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //732 padding zeros 42
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //733 padding zeros 43
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //734 padding zeros 44
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //735 padding zeros 45
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 

 //736 padding zeros 46
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //737 padding zeros 47
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //738 padding zeros 48
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //739 padding zeros 49
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //740 padding zeros 50
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //741 padding zeros 51
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //742 padding zeros 52
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //743 padding zeros 53
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //744 padding zeros 54
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //745 padding zeros 55
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 

 //746 padding zeros 56
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //747 padding zeros 57
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //748 padding zeros 58
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //749 padding zeros 59
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //750 padding zeros 60
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //751 padding zeros 61
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //752 padding zeros 62
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //753 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

 //754 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

 //755 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //756 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //757 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //758 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //759 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

 //760 padding zeros 60
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //761 padding zeros 61
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //762 padding zeros 62
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //763 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

 //764 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

 //765 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //766 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //767 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //768 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //769 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //770 padding zeros 60
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //771 padding zeros 61
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //772 padding zeros 62
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //773 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

 //774 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

 //775 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //776 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //777 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //778 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //779 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //780 padding zeros 60
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //781 padding zeros 61
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //782 padding zeros 62
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //783 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

 //784 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

 //785 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //786 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //787 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //788 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //789 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  //790 padding zeros 60
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //791 padding zeros 61
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //792 padding zeros 62
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //793 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

 //794 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

 //795 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //796 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //797 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //798 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //799 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //800 padding zeros  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 

 //801 padding zeros
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //802 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //803 padding zeros
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //804 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //805 padding zeros
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 

 //806 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //807 padding zeros
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //808 padding zeros
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //809 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //810 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 

 //811 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //812 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //813 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //814 padding zeros
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //815 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 

 //816 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //817 padding zeros
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //818 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //819 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //820 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //821 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //822 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //823 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //824 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //825 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 

 //826 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //827 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //828 padding zeros 38
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //829 padding zeros 39
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //830 padding zeros 40
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //831 padding zeros 41
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //832 padding zeros 42
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //833 padding zeros 43
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //834 padding zeros 44
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //835 padding zeros 45
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 

 //836 padding zeros 46
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //837 padding zeros 47
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //838 padding zeros 48
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //839 padding zeros 49
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //840 padding zeros 50
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //841 padding zeros 51
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //842 padding zeros 52
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //843 padding zeros 53
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //844 padding zeros 54
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //845 padding zeros 55
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 

 //846 padding zeros 56
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //847 padding zeros 57
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //848 padding zeros 58
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //849 padding zeros 59
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //850 padding zeros 60
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //851 padding zeros 61
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //852 padding zeros 62
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //853 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

 //854 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

 //855 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //856 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //857 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //858 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //859 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

 //860 padding zeros 60
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //861 padding zeros 61
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //862 padding zeros 62
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //863 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

 //864 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

 //865 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //866 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //867 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //868 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //869 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //870 padding zeros 60
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //871 padding zeros 61
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //872 padding zeros 62
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //873 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

 //874 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

 //875 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //876 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //877 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //878 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //879 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //880 padding zeros 60
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //881 padding zeros 61
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //882 padding zeros 62
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //883 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

 //884 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

 //885 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //886 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //887 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //888 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //889 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  //890 padding zeros 60
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //891 padding zeros 61
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //892 padding zeros 62
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //893 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

 //894 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

 //895 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //896 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //897 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //898 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //899 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  //900 padding zeros  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 

 //901 padding zeros
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //902 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //903 padding zeros
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //904 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //905 padding zeros
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 

 //906 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //907 padding zeros
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //908 padding zeros
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //909 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //910 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 

 //911 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //912 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //913 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //914 padding zeros
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //915 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 

 //916 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //917 padding zeros
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //918 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //919 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //920 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //921 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //922 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //923 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //924 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //925 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 

 //926 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //927 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //928 padding zeros 38
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //929 padding zeros 39
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //930 padding zeros 40
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //931 padding zeros 41
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //932 padding zeros 42
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //933 padding zeros 43
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //934 padding zeros 44
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //935 padding zeros 45
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 

 //936 padding zeros 46
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //937 padding zeros 47
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //938 padding zeros 48
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //939 padding zeros 49
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //940 padding zeros 50
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //941 padding zeros 51
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //942 padding zeros 52
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //943 padding zeros 53
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //944 padding zeros 54
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //945 padding zeros 55
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 

 //946 padding zeros 56
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //947 padding zeros 57
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //948 padding zeros 58
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //949 padding zeros 59
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //950 padding zeros 60
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //951 padding zeros 61
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //952 padding zeros 62
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //953 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

 //954 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

 //955 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //956 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //957 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //958 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //959 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

 //960 padding zeros 60
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //961 padding zeros 61
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //962 padding zeros 62
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //963 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

 //964 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

 //965 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //966 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //967 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //968 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //969 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //970 padding zeros 60
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //971 padding zeros 61
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //972 padding zeros 62
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //973 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

 //974 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

 //975 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //976 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //977 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //978 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //979 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //980 padding zeros 60
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //981 padding zeros 61
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //982 padding zeros 62
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //983 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

 //984 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

 //985 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //986 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //987 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //988 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //989 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  //990 padding zeros 60
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //991 padding zeros 61
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //992 padding zeros 62
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //993 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

 //994 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

 //995 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //996 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //997 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //998 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //999 padding zeros 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  //1000 padding zeros  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 

 //1001 padding zeros
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //1002 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //1003 padding zeros
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //1004 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //1005 padding zeros
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 

 //1006 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //1007 padding zeros
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //1008 padding zeros
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //1009 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //1010 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 

 //1011 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //1012 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //1013 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //1014 padding zeros
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //1015 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 

 //1016 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //1017 padding zeros
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //1018 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //1019 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //1020 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //1021 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //1022 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //1023 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
 //1024 padding zeros 
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// d - length of hash arrive 
//1: e0
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  
  #104166   tb_RxD   = 1;

//2: 00  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

// Key 
// 1: 61
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

// 2: 62  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
// 3: 63
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
//4: 64
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//5: 65
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
//6: 31
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
//7: 32
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
//8: 33
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//9: 34
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//10: 35
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//11: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//12: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//13: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//14: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//15: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//16: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//17: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//18: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//19: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//20: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//21: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//22: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//23: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//24: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//25: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//26: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//27: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//28: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//29: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//30: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//31: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//32: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//33: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//34: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//35: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//36: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//37: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//38: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//39: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
//40: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//41: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//42: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//43: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//44: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//45: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//46: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//47: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//48: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//49: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//50: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//51: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//52: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//53: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//54: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//55: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//56: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//57: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//58: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//59: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//60: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//61: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//62: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//63: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//64: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

// L
//40
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1; //"=1" to get L=64
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

// r 
//1: 05
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//2: 00  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//   keylen
//0a
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

// index padding  
//1: 40
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1; 

//2: 0d
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

// index index pad  
//01
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  //transmit
  #500000    button_tx  = 1;  
end

always begin
   #5  tb_clk = ~tb_clk; 
end

// Connect DUT to test bench
top DUT 
(
tb_clk  ,
tb_reset,
button_tx,
tb_RxD,
tb_done_M,
tb_done_d,
tb_done_K,
tb_done_L,
tb_done_r,
tb_done_keylen,
tb_done_padding,
tb_done_rx,
tb_TxD
);
  
endmodule
