///////////////////////////////////
// Verilog testbench
///////////////////////////////////
//last update: 26/11/2023

`timescale	1ns/1ps

module tb_top
(
);
  reg tb_clk, tb_reset;
  reg button_tx;
  reg [7:0] tb_RxD;
  wire tb_done_M;
  wire tb_done_d;
  wire  tb_done_K;
  wire tb_done_L;
  wire tb_done_r;
  wire tb_done_keylen;
  wire tb_done_padding;
  wire tb_done_rx;
  wire tb_done_MD6;
  wire tb_TxD;
  
initial begin
//  $display ("time\t\t  clk reset	 btn 	 rx 	 tx   ");
//  $monitor ("%8g\t\t%b   %b    %b	%b	%b", 
//	  $time, tb_clk, tb_reset, button_tx , tb_RxD , tb_TxD);	        	
  tb_clk             = 1; 
  tb_reset           = 1;
  button_tx 		 = 0;
  #700   tb_reset    = 0;
  
// message arrival
  #0	    tb_RxD   = 1;
  
  //1: 61
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 1; 
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //2: 62
  #104166   tb_RxD   = 0;  
  
  #104166   tb_RxD   = 0; 
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;

  #104166   tb_RxD   = 1;

  //3:	63  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //4: 00  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //5: 00  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //6: 00  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //7: 00  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //8: 00
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //9: 00
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //10: 00  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //11: 00  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //12: "55"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //13: "66"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //14: "77"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //15 "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //16: "22"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //17: "33" - 13  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //18: "44"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //19: "55"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //20: "66"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //21: "77"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //22: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //23: "22"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //24: "33"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //25: "44" - 14  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //26: "55"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //27: "66"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //28: "77"  
   #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //29: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //30 "22"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //31: "33"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //32: "44"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //33: "55" - 15  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //34: "66"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //35: "77"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //36: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //37: "22"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //38: "33"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //39: "44"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //40: "55"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //41: "66" - 16  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //42: "77"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //43: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //44: "22"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //45: "33"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //46: "44"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //47: "55"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //48: "66"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //49: "77" - 17  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //50: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //51: "22"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //52: "33"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //53: "44"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //54: "55"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //55: "66"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //56: "77"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //57: "11" - 21
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //58: "22"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //59: "33"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //60: "44"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //61: "55"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //62: "66"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //63: "77"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //64: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //65: "22" - 22
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //66: "33"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //67: "44"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //68: "55"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //69: "66"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //70: "77"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //71: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //72: "22"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //73: "33" - 23  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //74: "44"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //75: "55"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //76: "66"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //77: "77"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //78: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //79: "22" 
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //80: "33"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //81: "44" - 24 
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //82: "55"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //83: "66"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //84: "77"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //85: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //86: "22"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //87: "33"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //88: "44"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //89: "55" - 25  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //90: "66"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //91: "77"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //92: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //93: "22"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //94: "33"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //95: "44"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //96: "55"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //97: "66" - 26  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //98: "77"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //99: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //100: "22"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //101: "33"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //102: "44"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //103: "55"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //104: "66"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //105: "77" - 27  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //106: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //107: "22" 
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //108: "33"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //109: "44"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //110: "55"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //111: "66"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //112: "77"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //113: "11" - 31
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //114: "22"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //115: "33"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //116: "44"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //117: "55"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //118: "66"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //119: "77"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //120: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //121: "22" - 32
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //122: "33"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //123: "44"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //124: "55"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //125: "66"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //126: "77"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //127: "11" 
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //128: "22"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //129: "33" - 33 
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //130: "44"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //131: "55"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //132: "66"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //133: "77"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //134: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //135: "22"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //136: "33"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //137: "44" - 34  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //138: "55"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //139: "66"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //140: "77"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //141: "11" - 11
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //142: "22"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //143: "33"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //144: "44"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //145: "55" - 35  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //146: "66"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //147: "77"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //148: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //149: "22"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //150: "33"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //151: "44"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //152: "55"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //153: "66" - 36  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //154: "77"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //155: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //156: "22"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //157: "33"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //158: "44"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //159: "55"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //160: "66"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //161: "77" - 37  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //162: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //163: "22"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //164: "33"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //165: "44"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //166: "55"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //167: "66"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //168: "77"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //169: "11" - 41
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //170: "22"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //171: "33"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //172: "44"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //173: "55"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //174: "66"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //175: "77"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //176: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //177: "22" - 42
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //178: "33"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //179: "44"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //180: "55"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //181: "66"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //182: "77"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //183: "11" 
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //184: "22"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //185: "33" - 43  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //186: "44"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //187: "55"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //188: "66"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //189: "77"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //190: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //191: "22"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //192: "33"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //193: "44" - 44  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //194: "55"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //195: "66"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //196: "77"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //197: "11" - 11
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //198: "22"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //199: "33"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //200: "44"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //201: "55" - 45
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //202: "66"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //203: "77"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //204: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //205: "22" 
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //206: "33"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //207: "44"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //208: "55"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //209: "66"  - 46 
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //210: "77"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //211: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //212: "22"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //213: "33"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //214: "44"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //215: "55"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //216: "66"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //217: "77" - 47  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //218: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //219: "22" 
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //220: "33"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //221: "44"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //222: "55"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //223: "66"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //224: "77"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //225: "11" - 51
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //226: "22"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //227: "33"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //228: "44"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //229: "55"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //230: "66"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //231: "77"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //232: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //233: "22" - 52
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //234: "33"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //235: "44"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //236: "55"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //237: "66"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //238: "77"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //239: "11" - 11
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //240: "22"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //241: "33" - 53  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //242: "44"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //243: "55"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //244: "66"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //245: "77"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //246: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //247: "22"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //248: "33"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //249:"44" - 54  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //250: "55"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //251: "66"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //252: "77"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //253: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //254: "22"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //255: "33"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //256: "44"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //257: "55" - 55  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //258: "66"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //259: "77"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //260: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //261: "22" 
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //262: "33"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //263: "44"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //264: "55"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //265: "66" - 56 
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //266: "77"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //267: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //268: "22"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //269: "33"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //270: "44"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //271: "55"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //272: "66"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //273: "77" - 57  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //274: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //275: "22"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //276: "33"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //277: "44"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //278: "55"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //279: "66"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //280: "77"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //281: "11" - 61
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //282: "22"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //283: "33"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //284: "44"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //285: "55"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //286: "66"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //287: "77"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //288: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //289: "22" - 62
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //290: "33"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //291: "44"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //292: "55"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //293: "66"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //294: "77"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //295: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //296: "22"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //297: "33" - 63  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //298: "44"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //299: "55"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //300: "66"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //301: "77"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //302: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //303: "22"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //304: "33"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //305: "44" - 64  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //306: "55"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //307 :"66"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //308: "77"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //309: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //310: "22"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //311: "33"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //312: "44"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //313: "55" - 65  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //314: "66"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //315: "77"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //316: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //317: "22"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //318: "33"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //319: "44"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //320: "55"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //321: "66" - 66  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //322: "77"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //323: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //324: "22"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //325: "33"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //326: "44"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //327: "55"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //328: "66"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //329: "77" - 67  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //330: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //331: "22"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //332: "33"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //333: "44"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //334: "55"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //335: "66"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //336: "77"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //337: "11" - 71
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //338: "22"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //339: "33"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //340: "44"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //341: "55"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //342: "66"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //343: "77"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //344: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //345: "22" - 72
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //346: "33"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //347: "44"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //348: "55"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //349: "66"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //350: "77"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //351: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //352: "22"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //353: "33" - 73  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //354: "44"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //355: "55"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //356: "66"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //357: "77"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //358: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //359: "22"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //360: "33"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //361: "44" - 74  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //362: "55"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //363: "66"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //364: "77"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //365: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //366: "22"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //367: "33"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //368: "44"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //369: "55" - 75  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //370: "66"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //371: "77"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //372: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //373: "22" - 12
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //374: "33"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //375: "44"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //376: "55"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //377: "66" - 76  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //378: "77"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //379: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //380: "22"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //381: "33"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //382: "44"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //383: "55"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //384: "66"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //385: "77" - 77  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //386: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //387: "22"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //388: "33"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //389: "44"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //390: "55"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //391: "66"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //392: "77"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //393: "11" - 81
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //394: "22"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //395: "33"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //396: "44"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //397: "55"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //398: "66"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //399: "77"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //400: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //401: "22" - 82
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //402: "33"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //403: "44"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //404: "55"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //405: "66"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //406: "77"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //407: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //408: "22"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //409: "33" - 83  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //410: "44"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //411: "55"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //412: "66"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //413: "77"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //414: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //415: "22"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //416: "33"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //417: "44" - 84  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //418: "55"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //419: "66"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //420: "77"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //421: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //422: "22"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //423: "33"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //424: "44"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //425: "55" - 85  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //426: "66"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //427: "77"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //428: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //429: "22"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //430: "33"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //431: "44"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //432: "55"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //433: "66" - 86  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //434: "77"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //435: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //436: "22"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //437: "33"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //438: "44"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //439: "55"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //440: "66"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //441: "77" - 87  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //442: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //443: "22"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //444: "33"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //445: "44"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //446: "55"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //447: "66"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //448: "77"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
   //449: "11" - 91
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //450: "22"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //451: "33"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //452: "44"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //453: "55"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //454: "66"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //455: "77"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //456: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //457: "22" - 92
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //458: "33"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //459: "44"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //460: "55"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //461: "66"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //462: "77"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //463: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //464: "22"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //465: "33" - 93  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //466: "44"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //467: "55"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //468: "66"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //469: "77"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //470: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //471: "22"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //472: "33"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //473: "44" - 94  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //474: "55"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //475: "66"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //476: "77"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //477: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //478: "22"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //479: "33"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //480: "44"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //481: "55" - 95  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //482: "66"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //483: "77"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //484: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //485: "22"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //486: "33"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //487: "44"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //488: "55"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //489: "66" - 96  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //490: "77"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //491: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //492: "22"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //493: "33"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //494: "44"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //495: "55"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //496: "66"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //497: "77" - 97  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //498: "11"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
  //499: "22"
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //500: "33"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //501: "44"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //502: "55"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //503: "66"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //504: "77"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
 
  //505: "11" - 101
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //506: 00
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //507: 00  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //508: 00  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //509: "00"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //510: "00"  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //511: 00  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

  //512: 00
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// d - length of hash arrive 
//1: 00
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//2: 01  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

// Key 
// 1: 00
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

// 2: 00  
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
// 3: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
//4: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//5: 00
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
//6: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
//7: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  
//8: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//9: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//10: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//11: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//12: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//13: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//14: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//15: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//16: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//17: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//18: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//19: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//20: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//21: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//22: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//23: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//24: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//25: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//26: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//27: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//28: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//29: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//30: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//31: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//32: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//33: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//34: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//35: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//36: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//37: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//38: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//39: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
//40: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//41: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//42: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//43: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//44: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//45: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//46: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//47: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//48: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//49: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//50: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//51: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//52: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//53: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//54: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//55: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//56: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//57: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//58: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//59: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//60: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//61: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//62: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//63: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//64: 00
  #104166   tb_RxD   = 0; 
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

// L
//40
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1; //"=1" to get L=64
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

// r 
//1: 05
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//2: 00  
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

//   keylen
//00
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

// index padding  
//1: e8
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  
  #104166   tb_RxD   = 1; 

//2: 0f
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 1;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;

// index index pad  
//00
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  #104166   tb_RxD   = 0;
  
  #104166   tb_RxD   = 1;
  //transmit
  #500000    button_tx  = 1;  
end

always begin
   #5  tb_clk = ~tb_clk; 
end

// Connect DUT to test bench
top DUT 
(
tb_clk  ,
tb_reset,
button_tx,
tb_RxD,
tb_done_M,
tb_done_d,
tb_done_K,
tb_done_L,
tb_done_r,
tb_done_keylen,
tb_done_padding,
tb_done_rx,
tb_done_MD6,
tb_TxD
);
  
endmodule
